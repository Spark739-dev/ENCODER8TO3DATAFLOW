library verilog;
use verilog.vl_types.all;
entity encoder8_vlg_vec_tst is
end encoder8_vlg_vec_tst;
