library verilog;
use verilog.vl_types.all;
entity encoder8_vlg_sample_tst is
    port(
        d0              : in     vl_logic;
        d1              : in     vl_logic;
        d2              : in     vl_logic;
        d3              : in     vl_logic;
        d4              : in     vl_logic;
        d5              : in     vl_logic;
        d6              : in     vl_logic;
        d7              : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end encoder8_vlg_sample_tst;
