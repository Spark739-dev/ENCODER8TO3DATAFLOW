library verilog;
use verilog.vl_types.all;
entity encoder8_vlg_check_tst is
    port(
        a0              : in     vl_logic;
        a1              : in     vl_logic;
        a2              : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end encoder8_vlg_check_tst;
